module voltage_to_temp(input wire clk,
                       input wire [11:0] voltage,
                       output reg [10:0] temp_c_signed,
                       output reg [11:0] temp_f_signed);

always @(posedge clk)
    if (voltage < 12'ha6e)  temp_c_signed[10] <= 1;   //c temp is negative
    else                    temp_c_signed[10] <= 0;   //c temp is positive

always @(posedge clk)
    if (voltage < 12'd2370) temp_f_signed[11] <= 1;   //f temp is negative
    else                    temp_f_signed[11] <= 0;   //f temp is positive

always @(posedge clk)
    if      (voltage < 12'h7d0) temp_c_signed[9:0] <= 10'd0;
    else if (voltage < 12'h7D9)	temp_c_signed[9:0] <=	10'd400;
    else if (voltage < 12'h7E4)	temp_c_signed[9:0] <=	10'd394;
    else if (voltage < 12'h7ED)	temp_c_signed[9:0] <=	10'd388;
    else if (voltage < 12'h7F8)	temp_c_signed[9:0] <=	10'd382;
    else if (voltage < 12'h802)	temp_c_signed[9:0] <=	10'd376;
    else if (voltage < 12'h80C)	temp_c_signed[9:0] <=	10'd370;
    else if (voltage < 12'h816)	temp_c_signed[9:0] <=	10'd364;
    else if (voltage < 12'h820)	temp_c_signed[9:0] <=	10'd358;
    else if (voltage < 12'h82A)	temp_c_signed[9:0] <=	10'd352;
    else if (voltage < 12'h834)	temp_c_signed[9:0] <=	10'd346;
    else if (voltage < 12'h83E)	temp_c_signed[9:0] <=	10'd340;
    else if (voltage < 12'h848)	temp_c_signed[9:0] <=	10'd334;
    else if (voltage < 12'h852)	temp_c_signed[9:0] <=	10'd328;
    else if (voltage < 12'h85C)	temp_c_signed[9:0] <=	10'd322;
    else if (voltage < 12'h866)	temp_c_signed[9:0] <=	10'd316;
    else if (voltage < 12'h870)	temp_c_signed[9:0] <=	10'd310;
    else if (voltage < 12'h87A)	temp_c_signed[9:0] <=	10'd304;
    else if (voltage < 12'h884)	temp_c_signed[9:0] <=	10'd298;
    else if (voltage < 12'h88E)	temp_c_signed[9:0] <=	10'd292;
    else if (voltage < 12'h898)	temp_c_signed[9:0] <=	10'd286;
    else if (voltage < 12'h8A2)	temp_c_signed[9:0] <=	10'd280;
    else if (voltage < 12'h8AC)	temp_c_signed[9:0] <=	10'd274;
    else if (voltage < 12'h8B6)	temp_c_signed[9:0] <=	10'd268;
    else if (voltage < 12'h8C0)	temp_c_signed[9:0] <=	10'd262;
    else if (voltage < 12'h8CA)	temp_c_signed[9:0] <=	10'd256;
    else if (voltage < 12'h8D4)	temp_c_signed[9:0] <=	10'd250;
    else if (voltage < 12'h8DE)	temp_c_signed[9:0] <=	10'd244;
    else if (voltage < 12'h8E8)	temp_c_signed[9:0] <=	10'd238;
    else if (voltage < 12'h8F2)	temp_c_signed[9:0] <=	10'd232;
    else if (voltage < 12'h8FC)	temp_c_signed[9:0] <=	10'd226;
    else if (voltage < 12'h906)	temp_c_signed[9:0] <=	10'd220;
    else if (voltage < 12'h910)	temp_c_signed[9:0] <=	10'd214;
    else if (voltage < 12'h91A)	temp_c_signed[9:0] <=	10'd208;
    else if (voltage < 12'h924)	temp_c_signed[9:0] <=	10'd202;
    else if (voltage < 12'h92E)	temp_c_signed[9:0] <=	10'd196;
    else if (voltage < 12'h938)	temp_c_signed[9:0] <=	10'd190;
    else if (voltage < 12'h942)	temp_c_signed[9:0] <=	10'd184;
    else if (voltage < 12'h94C)	temp_c_signed[9:0] <=	10'd178;
    else if (voltage < 12'h956)	temp_c_signed[9:0] <=	10'd172;
    else if (voltage < 12'h960)	temp_c_signed[9:0] <=	10'd166;
    else if (voltage < 12'h96A)	temp_c_signed[9:0] <=	10'd160;
    else if (voltage < 12'h974)	temp_c_signed[9:0] <=	10'd154;
    else if (voltage < 12'h97E)	temp_c_signed[9:0] <=	10'd148;
    else if (voltage < 12'h988)	temp_c_signed[9:0] <=	10'd142;
    else if (voltage < 12'h992)	temp_c_signed[9:0] <=	10'd136;
    else if (voltage < 12'h99C)	temp_c_signed[9:0] <=	10'd130;
    else if (voltage < 12'h9A6)	temp_c_signed[9:0] <=	10'd124;
    else if (voltage < 12'h9B0)	temp_c_signed[9:0] <=	10'd118;
    else if (voltage < 12'h9BA)	temp_c_signed[9:0] <=	10'd112;
    else if (voltage < 12'h9C4)	temp_c_signed[9:0] <=	10'd106;
    else if (voltage < 12'h9CE)	temp_c_signed[9:0] <=	10'd100;
    else if (voltage < 12'h9D8)	temp_c_signed[9:0] <=	10'd94;
    else if (voltage < 12'h9E2)	temp_c_signed[9:0] <=	10'd88;
    else if (voltage < 12'h9EC)	temp_c_signed[9:0] <=	10'd82;
    else if (voltage < 12'h9F6)	temp_c_signed[9:0] <=	10'd76;
    else if (voltage < 12'hA00)	temp_c_signed[9:0] <=	10'd70;
    else if (voltage < 12'hA0A)	temp_c_signed[9:0] <=	10'd64;
    else if (voltage < 12'hA14)	temp_c_signed[9:0] <=	10'd58;
    else if (voltage < 12'hA1E)	temp_c_signed[9:0] <=	10'd52;
    else if (voltage < 12'hA28)	temp_c_signed[9:0] <=	10'd46;
    else if (voltage < 12'hA32)	temp_c_signed[9:0] <=	10'd40;
    else if (voltage < 12'hA3C)	temp_c_signed[9:0] <=	10'd34;
    else if (voltage < 12'hA46)	temp_c_signed[9:0] <=	10'd28;
    else if (voltage < 12'hA50)	temp_c_signed[9:0] <=	10'd22;
    else if (voltage < 12'hA5A)	temp_c_signed[9:0] <=	10'd16;
    else if (voltage < 12'hA64)	temp_c_signed[9:0] <=	10'd10;
    else if (voltage < 12'hA6E)	temp_c_signed[9:0] <=	10'd4;
    else if (voltage < 12'hA78)	temp_c_signed[9:0] <=	10'd2;
    else if (voltage < 12'hA82)	temp_c_signed[9:0] <=	10'd8;
    else if (voltage < 12'hA8C)	temp_c_signed[9:0] <=	10'd14;
    else if (voltage < 12'hA96)	temp_c_signed[9:0] <=	10'd20;
    else if (voltage < 12'hAA0)	temp_c_signed[9:0] <=	10'd26;
    else if (voltage < 12'hAAA)	temp_c_signed[9:0] <=	10'd32;
    else if (voltage < 12'hAB4)	temp_c_signed[9:0] <=	10'd38;
    else if (voltage < 12'hABD)	temp_c_signed[9:0] <=	10'd44;
    else if (voltage < 12'hAC8)	temp_c_signed[9:0] <=	10'd50;
    else if (voltage < 12'hAD1)	temp_c_signed[9:0] <=	10'd56;
    else if (voltage < 12'hADB)	temp_c_signed[9:0] <=	10'd62;
    else if (voltage < 12'hAE5)	temp_c_signed[9:0] <=	10'd68;
    else if (voltage < 12'hAEF)	temp_c_signed[9:0] <=	10'd74;
    else if (voltage < 12'hAF9)	temp_c_signed[9:0] <=	10'd80;
    else if (voltage < 12'hB03)	temp_c_signed[9:0] <=	10'd86;
    else if (voltage < 12'hB0D)	temp_c_signed[9:0] <=	10'd92;
    else if (voltage < 12'hB17)	temp_c_signed[9:0] <=	10'd98;
    else if (voltage < 12'hB21)	temp_c_signed[9:0] <=	10'd104;
    else if (voltage < 12'hB2B)	temp_c_signed[9:0] <=	10'd110;
    else if (voltage < 12'hB35)	temp_c_signed[9:0] <=	10'd116;
    else if (voltage < 12'hB3F)	temp_c_signed[9:0] <=	10'd122;
    else if (voltage < 12'hB49)	temp_c_signed[9:0] <=	10'd128;
    else if (voltage < 12'hB53)	temp_c_signed[9:0] <=	10'd134;
    else if (voltage < 12'hB5D)	temp_c_signed[9:0] <=	10'd140;
    else if (voltage < 12'hB67)	temp_c_signed[9:0] <=	10'd146;
    else if (voltage < 12'hB71)	temp_c_signed[9:0] <=	10'd152;
    else if (voltage < 12'hB7B)	temp_c_signed[9:0] <=	10'd158;
    else if (voltage < 12'hB85)	temp_c_signed[9:0] <=	10'd164;
    else if (voltage < 12'hB8F)	temp_c_signed[9:0] <=	10'd170;
    else if (voltage < 12'hB99)	temp_c_signed[9:0] <=	10'd176;
    else if (voltage < 12'hBA3)	temp_c_signed[9:0] <=	10'd182;
    else if (voltage < 12'hBAD)	temp_c_signed[9:0] <=	10'd188;
    else if (voltage < 12'hBB7)	temp_c_signed[9:0] <=	10'd194;
    else if (voltage < 12'hBC1)	temp_c_signed[9:0] <=	10'd200;
    else if (voltage < 12'hBCB)	temp_c_signed[9:0] <=	10'd206;
    else if (voltage < 12'hBD5)	temp_c_signed[9:0] <=	10'd212;
    else if (voltage < 12'hBDF)	temp_c_signed[9:0] <=	10'd218;
    else if (voltage < 12'hBE9)	temp_c_signed[9:0] <=	10'd224;
    else if (voltage < 12'hBF3)	temp_c_signed[9:0] <=	10'd230;
    else if (voltage < 12'hBFD)	temp_c_signed[9:0] <=	10'd236;
    else if (voltage < 12'hC07)	temp_c_signed[9:0] <=	10'd242;
    else if (voltage < 12'hC11)	temp_c_signed[9:0] <=	10'd248;
    else if (voltage < 12'hC1B)	temp_c_signed[9:0] <=	10'd254;
    else if (voltage < 12'hC25)	temp_c_signed[9:0] <=	10'd260;
    else if (voltage < 12'hC2F)	temp_c_signed[9:0] <=	10'd266;
    else if (voltage < 12'hC39)	temp_c_signed[9:0] <=	10'd272;
    else if (voltage < 12'hC43)	temp_c_signed[9:0] <=	10'd278;
    else if (voltage < 12'hC4D)	temp_c_signed[9:0] <=	10'd284;
    else if (voltage < 12'hC57)	temp_c_signed[9:0] <=	10'd290;
    else if (voltage < 12'hC61)	temp_c_signed[9:0] <=	10'd296;
    else if (voltage < 12'hC6B)	temp_c_signed[9:0] <=	10'd302;
    else if (voltage < 12'hC75)	temp_c_signed[9:0] <=	10'd308;
    else if (voltage < 12'hC7F)	temp_c_signed[9:0] <=	10'd314;
    else if (voltage < 12'hC89)	temp_c_signed[9:0] <=	10'd320;
    else if (voltage < 12'hC93)	temp_c_signed[9:0] <=	10'd326;
    else if (voltage < 12'hC9D)	temp_c_signed[9:0] <=	10'd332;
    else if (voltage < 12'hCA7)	temp_c_signed[9:0] <=	10'd338;
    else if (voltage < 12'hCB1)	temp_c_signed[9:0] <=	10'd344;
    else if (voltage < 12'hCBB)	temp_c_signed[9:0] <=	10'd350;
    else if (voltage < 12'hCC5)	temp_c_signed[9:0] <=	10'd356;
    else if (voltage < 12'hCCF)	temp_c_signed[9:0] <=	10'd362;
    else if (voltage < 12'hCD9)	temp_c_signed[9:0] <=	10'd368;
    else if (voltage < 12'hCE3)	temp_c_signed[9:0] <=	10'd374;
    else if (voltage < 12'hCED)	temp_c_signed[9:0] <=	10'd380;
    else if (voltage < 12'hCF7)	temp_c_signed[9:0] <=	10'd386;
    else if (voltage < 12'hD01)	temp_c_signed[9:0] <=	10'd392;
    else if (voltage < 12'hD0B)	temp_c_signed[9:0] <=	10'd398;
    else if (voltage < 12'hD15)	temp_c_signed[9:0] <=	10'd404;
    else if (voltage < 12'hD1F)	temp_c_signed[9:0] <=	10'd410;
    else if (voltage < 12'hD29)	temp_c_signed[9:0] <=	10'd416;
    else if (voltage < 12'hD33)	temp_c_signed[9:0] <=	10'd422;
    else if (voltage < 12'hD3D)	temp_c_signed[9:0] <=	10'd428;
    else if (voltage < 12'hD47)	temp_c_signed[9:0] <=	10'd434;
    else if (voltage < 12'hD51)	temp_c_signed[9:0] <=	10'd440;
    else if (voltage < 12'hD5B)	temp_c_signed[9:0] <=	10'd446;
    else if (voltage < 12'hD65)	temp_c_signed[9:0] <=	10'd452;
    else if (voltage < 12'hD6F)	temp_c_signed[9:0] <=	10'd458;
    else if (voltage < 12'hD79)	temp_c_signed[9:0] <=	10'd464;
    else if (voltage < 12'hD83)	temp_c_signed[9:0] <=	10'd470;
    else if (voltage < 12'hD8D)	temp_c_signed[9:0] <=	10'd476;
    else if (voltage < 12'hD97)	temp_c_signed[9:0] <=	10'd482;
    else if (voltage < 12'hDA1)	temp_c_signed[9:0] <=	10'd488;
    else if (voltage < 12'hDAB)	temp_c_signed[9:0] <=	10'd494;
    else if (voltage < 12'hDB5)	temp_c_signed[9:0] <=	10'd500;
    else if (voltage < 12'hDBF)	temp_c_signed[9:0] <=	10'd506;
    else if (voltage < 12'hDC9)	temp_c_signed[9:0] <=	10'd512;
    else if (voltage < 12'hDD3)	temp_c_signed[9:0] <=	10'd518;
    else if (voltage < 12'hDDD)	temp_c_signed[9:0] <=	10'd524;
    else if (voltage < 12'hDE7)	temp_c_signed[9:0] <=	10'd530;
    else if (voltage < 12'hDF1)	temp_c_signed[9:0] <=	10'd536;
    else if (voltage < 12'hDFB)	temp_c_signed[9:0] <=	10'd542;
    else if (voltage < 12'hE05)	temp_c_signed[9:0] <=	10'd548;
    else if (voltage < 12'hE0F)	temp_c_signed[9:0] <=	10'd554;
    else if (voltage < 12'hE19)	temp_c_signed[9:0] <=	10'd560;
    else if (voltage < 12'hE23)	temp_c_signed[9:0] <=	10'd566;
    else if (voltage < 12'hE2D)	temp_c_signed[9:0] <=	10'd572;
    else if (voltage < 12'hE37)	temp_c_signed[9:0] <=	10'd578;
    else if (voltage < 12'hE41)	temp_c_signed[9:0] <=	10'd584;
    else if (voltage < 12'hE4B)	temp_c_signed[9:0] <=	10'd590;
    else if (voltage < 12'hE55)	temp_c_signed[9:0] <=	10'd596;
    else if (voltage < 12'hE5F)	temp_c_signed[9:0] <=	10'd602;
    else if (voltage < 12'hE69)	temp_c_signed[9:0] <=	10'd608;
    else if (voltage < 12'hE73)	temp_c_signed[9:0] <=	10'd614;
    else if (voltage < 12'hE7D)	temp_c_signed[9:0] <=	10'd620;
    else if (voltage < 12'hE87)	temp_c_signed[9:0] <=	10'd626;
    else if (voltage < 12'hE91)	temp_c_signed[9:0] <=	10'd632;
    else if (voltage < 12'hE9B)	temp_c_signed[9:0] <=	10'd638;
    else if (voltage < 12'hEA5)	temp_c_signed[9:0] <=	10'd644;
    else if (voltage < 12'hEAF)	temp_c_signed[9:0] <=	10'd650;
    else if (voltage < 12'hEB9)	temp_c_signed[9:0] <=	10'd656;
    else if (voltage < 12'hEC3)	temp_c_signed[9:0] <=	10'd662;
    else if (voltage < 12'hECD)	temp_c_signed[9:0] <=	10'd668;
    else if (voltage < 12'hED7)	temp_c_signed[9:0] <=	10'd674;
    else if (voltage < 12'hEE1)	temp_c_signed[9:0] <=	10'd680;
    else if (voltage < 12'hEEB)	temp_c_signed[9:0] <=	10'd686;
    else if (voltage < 12'hEF5)	temp_c_signed[9:0] <=	10'd692;
    else if (voltage < 12'hEFF)	temp_c_signed[9:0] <=	10'd698;
    else if (voltage < 12'hF09)	temp_c_signed[9:0] <=	10'd704;
    else if (voltage < 12'hF13)	temp_c_signed[9:0] <=	10'd710;
    else if (voltage < 12'hF1D)	temp_c_signed[9:0] <=	10'd716;
    else if (voltage < 12'hF27)	temp_c_signed[9:0] <=	10'd722;
    else if (voltage < 12'hF31)	temp_c_signed[9:0] <=	10'd728;
    else if (voltage < 12'hF3B)	temp_c_signed[9:0] <=	10'd734;
    else if (voltage < 12'hF45)	temp_c_signed[9:0] <=	10'd740;
    else if (voltage < 12'hF4F)	temp_c_signed[9:0] <=	10'd746;
    else if (voltage < 12'hF59)	temp_c_signed[9:0] <=	10'd752;
    else if (voltage < 12'hF63)	temp_c_signed[9:0] <=	10'd758;
    else if (voltage < 12'hF6D)	temp_c_signed[9:0] <=	10'd764;
    else if (voltage < 12'hF77)	temp_c_signed[9:0] <=	10'd770;
    else if (voltage < 12'hF81)	temp_c_signed[9:0] <=	10'd776;
    else if (voltage < 12'hF8B)	temp_c_signed[9:0] <=	10'd782;
    else if (voltage < 12'hF95)	temp_c_signed[9:0] <=	10'd788;
    else if (voltage < 12'hF9F)	temp_c_signed[9:0] <=	10'd794;
    else                        temp_c_signed[9:0] <=	10'd0;

always @(posedge clk)
    if (voltage < 12'h7d0)      temp_f_signed[10:0] <= 10'd0;
    else if (voltage < 12'h7E4)	temp_f_signed[10:0] <=	10'd400;
    else if (voltage < 12'h7ED)	temp_f_signed[10:0] <=	10'd389;
    else if (voltage < 12'h7F8)	temp_f_signed[10:0] <=	10'd378;
    else if (voltage < 12'h802)	temp_f_signed[10:0] <=	10'd368;
    else if (voltage < 12'h80C)	temp_f_signed[10:0] <=	10'd357;
    else if (voltage < 12'h816)	temp_f_signed[10:0] <=	10'd346;
    else if (voltage < 12'h820)	temp_f_signed[10:0] <=	10'd335;
    else if (voltage < 12'h82A)	temp_f_signed[10:0] <=	10'd324;
    else if (voltage < 12'h834)	temp_f_signed[10:0] <=	10'd314;
    else if (voltage < 12'h83E)	temp_f_signed[10:0] <=	10'd303;
    else if (voltage < 12'h848)	temp_f_signed[10:0] <=	10'd292;
    else if (voltage < 12'h852)	temp_f_signed[10:0] <=	10'd281;
    else if (voltage < 12'h85C)	temp_f_signed[10:0] <=	10'd270;
    else if (voltage < 12'h866)	temp_f_signed[10:0] <=	10'd260;
    else if (voltage < 12'h870)	temp_f_signed[10:0] <=	10'd249;
    else if (voltage < 12'h87A)	temp_f_signed[10:0] <=	10'd238;
    else if (voltage < 12'h884)	temp_f_signed[10:0] <=	10'd227;
    else if (voltage < 12'h88E)	temp_f_signed[10:0] <=	10'd216;
    else if (voltage < 12'h898)	temp_f_signed[10:0] <=	10'd206;
    else if (voltage < 12'h8A2)	temp_f_signed[10:0] <=	10'd195;
    else if (voltage < 12'h8AC)	temp_f_signed[10:0] <=	10'd184;
    else if (voltage < 12'h8B6)	temp_f_signed[10:0] <=	10'd173;
    else if (voltage < 12'h8C0)	temp_f_signed[10:0] <=	10'd162;
    else if (voltage < 12'h8CA)	temp_f_signed[10:0] <=	10'd152;
    else if (voltage < 12'h8D4)	temp_f_signed[10:0] <=	10'd141;
    else if (voltage < 12'h8DE)	temp_f_signed[10:0] <=	10'd130;
    else if (voltage < 12'h8E8)	temp_f_signed[10:0] <=	10'd119;
    else if (voltage < 12'h8F2)	temp_f_signed[10:0] <=	10'd108;
    else if (voltage < 12'h8FC)	temp_f_signed[10:0] <=	10'd98;
    else if (voltage < 12'h906)	temp_f_signed[10:0] <=	10'd87;
    else if (voltage < 12'h910)	temp_f_signed[10:0] <=	10'd76;
    else if (voltage < 12'h91A)	temp_f_signed[10:0] <=	10'd65;
    else if (voltage < 12'h924)	temp_f_signed[10:0] <=	10'd54;
    else if (voltage < 12'h92E)	temp_f_signed[10:0] <=	10'd44;
    else if (voltage < 12'h938)	temp_f_signed[10:0] <=	10'd33;
    else if (voltage < 12'h942)	temp_f_signed[10:0] <=	10'd22;
    else if (voltage < 12'h94C)	temp_f_signed[10:0] <=	10'd11;
    else if (voltage < 12'h956)	temp_f_signed[10:0] <=	10'd0;
    else if (voltage < 12'h960)	temp_f_signed[10:0] <=	10'd10;
    else if (voltage < 12'h96A)	temp_f_signed[10:0] <=	10'd21;
    else if (voltage < 12'h974)	temp_f_signed[10:0] <=	10'd32;
    else if (voltage < 12'h97E)	temp_f_signed[10:0] <=	10'd43;
    else if (voltage < 12'h988)	temp_f_signed[10:0] <=	10'd54;
    else if (voltage < 12'h992)	temp_f_signed[10:0] <=	10'd64;
    else if (voltage < 12'h99C)	temp_f_signed[10:0] <=	10'd75;
    else if (voltage < 12'h9A6)	temp_f_signed[10:0] <=	10'd86;
    else if (voltage < 12'h9B0)	temp_f_signed[10:0] <=	10'd97;
    else if (voltage < 12'h9BA)	temp_f_signed[10:0] <=	10'd108;
    else if (voltage < 12'h9C4)	temp_f_signed[10:0] <=	10'd118;
    else if (voltage < 12'h9CE)	temp_f_signed[10:0] <=	10'd129;
    else if (voltage < 12'h9D8)	temp_f_signed[10:0] <=	10'd140;
    else if (voltage < 12'h9E2)	temp_f_signed[10:0] <=	10'd151;
    else if (voltage < 12'h9EC)	temp_f_signed[10:0] <=	10'd162;
    else if (voltage < 12'h9F6)	temp_f_signed[10:0] <=	10'd172;
    else if (voltage < 12'hA00)	temp_f_signed[10:0] <=	10'd183;
    else if (voltage < 12'hA0A)	temp_f_signed[10:0] <=	10'd194;
    else if (voltage < 12'hA14)	temp_f_signed[10:0] <=	10'd205;
    else if (voltage < 12'hA1E)	temp_f_signed[10:0] <=	10'd216;
    else if (voltage < 12'hA28)	temp_f_signed[10:0] <=	10'd226;
    else if (voltage < 12'hA32)	temp_f_signed[10:0] <=	10'd237;
    else if (voltage < 12'hA3C)	temp_f_signed[10:0] <=	10'd248;
    else if (voltage < 12'hA46)	temp_f_signed[10:0] <=	10'd259;
    else if (voltage < 12'hA50)	temp_f_signed[10:0] <=	10'd270;
    else if (voltage < 12'hA5A)	temp_f_signed[10:0] <=	10'd280;
    else if (voltage < 12'hA64)	temp_f_signed[10:0] <=	10'd291;
    else if (voltage < 12'hA6E)	temp_f_signed[10:0] <=	10'd302;
    else if (voltage < 12'hA78)	temp_f_signed[10:0] <=	10'd313;
    else if (voltage < 12'hA82)	temp_f_signed[10:0] <=	10'd324;
    else if (voltage < 12'hA8C)	temp_f_signed[10:0] <=	10'd334;
    else if (voltage < 12'hA96)	temp_f_signed[10:0] <=	10'd345;
    else if (voltage < 12'hAA0)	temp_f_signed[10:0] <=	10'd356;
    else if (voltage < 12'hAAA)	temp_f_signed[10:0] <=	10'd367;
    else if (voltage < 12'hAB4)	temp_f_signed[10:0] <=	10'd378;
    else if (voltage < 12'hABD)	temp_f_signed[10:0] <=	10'd388;
    else if (voltage < 12'hAC8)	temp_f_signed[10:0] <=	10'd399;
    else if (voltage < 12'hAD1)	temp_f_signed[10:0] <=	10'd410;
    else if (voltage < 12'hADB)	temp_f_signed[10:0] <=	10'd421;
    else if (voltage < 12'hAE5)	temp_f_signed[10:0] <=	10'd432;
    else if (voltage < 12'hAEF)	temp_f_signed[10:0] <=	10'd442;
    else if (voltage < 12'hAF9)	temp_f_signed[10:0] <=	10'd453;
    else if (voltage < 12'hB03)	temp_f_signed[10:0] <=	10'd464;
    else if (voltage < 12'hB0D)	temp_f_signed[10:0] <=	10'd475;
    else if (voltage < 12'hB17)	temp_f_signed[10:0] <=	10'd486;
    else if (voltage < 12'hB21)	temp_f_signed[10:0] <=	10'd496;
    else if (voltage < 12'hB2B)	temp_f_signed[10:0] <=	10'd507;
    else if (voltage < 12'hB35)	temp_f_signed[10:0] <=	10'd518;
    else if (voltage < 12'hB3F)	temp_f_signed[10:0] <=	10'd529;
    else if (voltage < 12'hB49)	temp_f_signed[10:0] <=	10'd540;
    else if (voltage < 12'hB53)	temp_f_signed[10:0] <=	10'd550;
    else if (voltage < 12'hB5D)	temp_f_signed[10:0] <=	10'd561;
    else if (voltage < 12'hB67)	temp_f_signed[10:0] <=	10'd572;
    else if (voltage < 12'hB71)	temp_f_signed[10:0] <=	10'd583;
    else if (voltage < 12'hB7B)	temp_f_signed[10:0] <=	10'd594;
    else if (voltage < 12'hB85)	temp_f_signed[10:0] <=	10'd604;
    else if (voltage < 12'hB8F)	temp_f_signed[10:0] <=	10'd615;
    else if (voltage < 12'hB99)	temp_f_signed[10:0] <=	10'd626;
    else if (voltage < 12'hBA3)	temp_f_signed[10:0] <=	10'd637;
    else if (voltage < 12'hBAD)	temp_f_signed[10:0] <=	10'd648;
    else if (voltage < 12'hBB7)	temp_f_signed[10:0] <=	10'd658;
    else if (voltage < 12'hBC1)	temp_f_signed[10:0] <=	10'd669;
    else if (voltage < 12'hBCB)	temp_f_signed[10:0] <=	10'd680;
    else if (voltage < 12'hBD5)	temp_f_signed[10:0] <=	10'd691;
    else if (voltage < 12'hBDF)	temp_f_signed[10:0] <=	10'd702;
    else if (voltage < 12'hBE9)	temp_f_signed[10:0] <=	10'd712;
    else if (voltage < 12'hBF3)	temp_f_signed[10:0] <=	10'd723;
    else if (voltage < 12'hBFD)	temp_f_signed[10:0] <=	10'd734;
    else if (voltage < 12'hC07)	temp_f_signed[10:0] <=	10'd745;
    else if (voltage < 12'hC11)	temp_f_signed[10:0] <=	10'd756;
    else if (voltage < 12'hC1B)	temp_f_signed[10:0] <=	10'd766;
    else if (voltage < 12'hC25)	temp_f_signed[10:0] <=	10'd777;
    else if (voltage < 12'hC2F)	temp_f_signed[10:0] <=	10'd788;
    else if (voltage < 12'hC39)	temp_f_signed[10:0] <=	10'd799;
    else if (voltage < 12'hC43)	temp_f_signed[10:0] <=	10'd810;
    else if (voltage < 12'hC4D)	temp_f_signed[10:0] <=	10'd820;
    else if (voltage < 12'hC57)	temp_f_signed[10:0] <=	10'd831;
    else if (voltage < 12'hC61)	temp_f_signed[10:0] <=	10'd842;
    else if (voltage < 12'hC6B)	temp_f_signed[10:0] <=	10'd853;
    else if (voltage < 12'hC75)	temp_f_signed[10:0] <=	10'd864;
    else if (voltage < 12'hC7F)	temp_f_signed[10:0] <=	10'd874;
    else if (voltage < 12'hC89)	temp_f_signed[10:0] <=	10'd885;
    else if (voltage < 12'hC93)	temp_f_signed[10:0] <=	10'd896;
    else if (voltage < 12'hC9D)	temp_f_signed[10:0] <=	10'd907;
    else if (voltage < 12'hCA7)	temp_f_signed[10:0] <=	10'd918;
    else if (voltage < 12'hCB1)	temp_f_signed[10:0] <=	10'd928;
    else if (voltage < 12'hCBB)	temp_f_signed[10:0] <=	10'd939;
    else if (voltage < 12'hCC5)	temp_f_signed[10:0] <=	10'd950;
    else if (voltage < 12'hCCF)	temp_f_signed[10:0] <=	10'd961;
    else if (voltage < 12'hCD9)	temp_f_signed[10:0] <=	10'd972;
    else if (voltage < 12'hCE3)	temp_f_signed[10:0] <=	10'd982;
    else if (voltage < 12'hCED)	temp_f_signed[10:0] <=	10'd993;
    else if (voltage < 12'hCF7)	temp_f_signed[10:0] <=	10'd1004;
    else if (voltage < 12'hD01)	temp_f_signed[10:0] <=	10'd1015;
    else if (voltage < 12'hD0B)	temp_f_signed[10:0] <=	10'd1026;
    else if (voltage < 12'hD15)	temp_f_signed[10:0] <=	10'd1036;
    else if (voltage < 12'hD1F)	temp_f_signed[10:0] <=	10'd1047;
    else if (voltage < 12'hD29)	temp_f_signed[10:0] <=	10'd1058;
    else if (voltage < 12'hD33)	temp_f_signed[10:0] <=	10'd1069;
    else if (voltage < 12'hD3D)	temp_f_signed[10:0] <=	10'd1080;
    else if (voltage < 12'hD47)	temp_f_signed[10:0] <=	10'd1090;
    else if (voltage < 12'hD51)	temp_f_signed[10:0] <=	10'd1101;
    else if (voltage < 12'hD5B)	temp_f_signed[10:0] <=	10'd1112;
    else if (voltage < 12'hD65)	temp_f_signed[10:0] <=	10'd1123;
    else if (voltage < 12'hD6F)	temp_f_signed[10:0] <=	10'd1134;
    else if (voltage < 12'hD79)	temp_f_signed[10:0] <=	10'd1144;
    else if (voltage < 12'hD83)	temp_f_signed[10:0] <=	10'd1155;
    else if (voltage < 12'hD8D)	temp_f_signed[10:0] <=	10'd1166;
    else if (voltage < 12'hD97)	temp_f_signed[10:0] <=	10'd1177;
    else if (voltage < 12'hDA1)	temp_f_signed[10:0] <=	10'd1188;
    else if (voltage < 12'hDAB)	temp_f_signed[10:0] <=	10'd1198;
    else if (voltage < 12'hDB5)	temp_f_signed[10:0] <=	10'd1209;
    else if (voltage < 12'hDBF)	temp_f_signed[10:0] <=	10'd1220;
    else if (voltage < 12'hDC9)	temp_f_signed[10:0] <=	10'd1231;
    else if (voltage < 12'hDD3)	temp_f_signed[10:0] <=	10'd1242;
    else if (voltage < 12'hDDD)	temp_f_signed[10:0] <=	10'd1252;
    else if (voltage < 12'hDE7)	temp_f_signed[10:0] <=	10'd1263;
    else if (voltage < 12'hDF1)	temp_f_signed[10:0] <=	10'd1274;
    else if (voltage < 12'hDFB)	temp_f_signed[10:0] <=	10'd1285;
    else if (voltage < 12'hE05)	temp_f_signed[10:0] <=	10'd1296;
    else if (voltage < 12'hE0F)	temp_f_signed[10:0] <=	10'd1306;
    else if (voltage < 12'hE19)	temp_f_signed[10:0] <=	10'd1317;
    else if (voltage < 12'hE23)	temp_f_signed[10:0] <=	10'd1328;
    else if (voltage < 12'hE2D)	temp_f_signed[10:0] <=	10'd1339;
    else if (voltage < 12'hE37)	temp_f_signed[10:0] <=	10'd1350;
    else if (voltage < 12'hE41)	temp_f_signed[10:0] <=	10'd1360;
    else if (voltage < 12'hE4B)	temp_f_signed[10:0] <=	10'd1371;
    else if (voltage < 12'hE55)	temp_f_signed[10:0] <=	10'd1382;
    else if (voltage < 12'hE5F)	temp_f_signed[10:0] <=	10'd1393;
    else if (voltage < 12'hE69)	temp_f_signed[10:0] <=	10'd1404;
    else if (voltage < 12'hE73)	temp_f_signed[10:0] <=	10'd1414;
    else if (voltage < 12'hE7D)	temp_f_signed[10:0] <=	10'd1425;
    else if (voltage < 12'hE87)	temp_f_signed[10:0] <=	10'd1436;
    else if (voltage < 12'hE91)	temp_f_signed[10:0] <=	10'd1447;
    else if (voltage < 12'hE9B)	temp_f_signed[10:0] <=	10'd1458;
    else if (voltage < 12'hEA5)	temp_f_signed[10:0] <=	10'd1468;
    else if (voltage < 12'hEAF)	temp_f_signed[10:0] <=	10'd1479;
    else if (voltage < 12'hEB9)	temp_f_signed[10:0] <=	10'd1490;
    else if (voltage < 12'hEC3)	temp_f_signed[10:0] <=	10'd1501;
    else if (voltage < 12'hECD)	temp_f_signed[10:0] <=	10'd1512;
    else if (voltage < 12'hED7)	temp_f_signed[10:0] <=	10'd1522;
    else if (voltage < 12'hEE1)	temp_f_signed[10:0] <=	10'd1533;
    else if (voltage < 12'hEEB)	temp_f_signed[10:0] <=	10'd1544;
    else if (voltage < 12'hEF5)	temp_f_signed[10:0] <=	10'd1555;
    else if (voltage < 12'hEFF)	temp_f_signed[10:0] <=	10'd1566;
    else if (voltage < 12'hF09)	temp_f_signed[10:0] <=	10'd1576;
    else if (voltage < 12'hF13)	temp_f_signed[10:0] <=	10'd1587;
    else if (voltage < 12'hF1D)	temp_f_signed[10:0] <=	10'd1598;
    else if (voltage < 12'hF27)	temp_f_signed[10:0] <=	10'd1609;
    else if (voltage < 12'hF31)	temp_f_signed[10:0] <=	10'd1620;
    else if (voltage < 12'hF3B)	temp_f_signed[10:0] <=	10'd1630;
    else if (voltage < 12'hF45)	temp_f_signed[10:0] <=	10'd1641;
    else if (voltage < 12'hF4F)	temp_f_signed[10:0] <=	10'd1652;
    else if (voltage < 12'hF59)	temp_f_signed[10:0] <=	10'd1663;
    else if (voltage < 12'hF63)	temp_f_signed[10:0] <=	10'd1674;
    else if (voltage < 12'hF6D)	temp_f_signed[10:0] <=	10'd1684;
    else if (voltage < 12'hF77)	temp_f_signed[10:0] <=	10'd1695;
    else if (voltage < 12'hF81)	temp_f_signed[10:0] <=	10'd1706;
    else if (voltage < 12'hF8B)	temp_f_signed[10:0] <=	10'd1717;
    else if (voltage < 12'hF95)	temp_f_signed[10:0] <=	10'd1728;
    else if (voltage < 12'hF9F)	temp_f_signed[10:0] <=	10'd1738;
    else                        temp_f_signed[10:0] <=   10'd0;

endmodule